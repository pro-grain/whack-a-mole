`timescale 1ns / 1ps

module timer(
    input clk,
    input rst_n,
    input load,
    input [3:0] load_tens_digit,
    input [3:0] load_ones_digit,
    output [3:0] tens_digit,
    output [3:0] ones_digit
    );
    
endmodule
