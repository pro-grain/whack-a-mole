`timescale 1ns / 1ps

module rand_gen(
    input clk,
    input rst_n,
    output [4:0] rand
    );
endmodule
