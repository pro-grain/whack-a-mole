`timescale 1ns / 1ps

module button(
    input clk,
    input rst_n,
    input raw_button,
    output button
    );
endmodule
