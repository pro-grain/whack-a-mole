`timescale 1ns / 1ps

module board_timer(
    input clk,
    input rst_n,
    input load,
    input [27:0] loadval,
    output time_trigger
    );
    
endmodule
