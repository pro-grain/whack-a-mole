`timescale 1ns / 1ps

module global_state(

    );
endmodule
